module shiftTest();

endmodule
