`include "alu.v"
`include "arithmetic.v"
`include "control_module.v"
`include "mux.v"
`include "doubleLeftShift.v"
`include "signExtendu.v"
`include "signExtends.v"
`include "regfile.v"
`include "datamemory.v"
`include "instrmemory.v"
module mips_cpu
(
  input clk
);
	wire[31:0] mem_read, alu_res, next_instruction_addr, instruction_addr, instruction_addr_plus4, 
				jumped_pc, extended_immediate, shifted_extended_immediate, b,
				normal_pc, pc_jump_addr, read_1, read_2, normal_write_data;
	wire[31:26] op;
	wire[25:21] rs;
	wire[25:0] jump_instruction_addr;
	wire[27:0] jump_instruction_addr_shifted;
	wire[20:16] rt;
	wire[15:11] rd;
	wire[10:6] shft;
	wire[5:0] func;
	wire[15:0] imm;
	wire[4:0] write_addr;
	wire[2:0] alu_op;
	wire reg_dest, alu_src, zero_flag, alu_op, write_enable, mem_write_enable, mem_read_enable, mem_to_reg, 
		 pc_src, jump_enable, bne_pc_override, pc_choose, jal_reg_override, normal_write_addr, overflow, carryout;
		 //carryout and overflow do nothing. We just need them for the ALU

	//Control Module
	cpu_control control_module(op, func, reg_dest, alu_src, mem_write_enable, mem_to_reg, pc_src, write_enable, mem_read_enable, alu_op, jump_enable, bne_pc_override, jal_reg_override); //checked

	//2:1 mux
	//ties pc_chooser mux directly to zero flag of ALU for use in BNE operations
	// input 0, input 1, choice, output
	mux #(2) bne_pc_override_mux(pc_src, zero_flag, bne_pc_override, pc_choose); //checked

	//PC register
	register32 PC(instruction_addr, next_instruction_addr, 1`b1, clk); //checked

	//PC incrementer
	bitwiseADD pc_incrementer(instruction_addr_plus4, overflow, instruction_addr, 32'd4, 1'b0); //checked

	//PC adder
	bitwiseADD pc_jumper(instruction_addr_plus_immediate, overflow, instruction_addr_plus4, shifted_extended_immediate, 1'b0); //checked

	//PC chooser
	mux #(32) pc_chooser(instruction_addr_plus4, instruction_addr_plus_immediate, pc_choose, normal_pc); //checked

	//PC Jumper
	mux #(32) jump_mux(normal_pc, pc_jump_addr, jump_enable, next_instruction_addr); //checked

	//Take address from instruction and shift left by 2
	doubleLeftShift jump_shifter(jump_instruction_addr, jump_instruction_addr_shifted, 1, clk); //checked

	//Concat shifted jump address with 4 most significant bits of PC+4
	//Stick the 4 most significant bits of PC+4 on to the shifted immediate from the instruction
	concatenator jump_add_concat(instruction_addr_plus4, jump_instruction_addr_shifted, clk, pc_jump_addr); //checked

	//instruction memory module
	#1
	instrmemory instruction_memory(instruction_addr, op, rs, rt, rd, shft, func, imm, jump_instruction_addr); //checked

	//instruction register destination mux
    //output, choice 1, choice 2, selector
	mux #(5) reg_dest_mux(rt, rd, reg_dest, normal_write_addr); //checked

	//mux to choose address to write to for jal op
	mux #(5) jal_reg_mux(normal_write_addr, 5'd31, jal_reg_override, write_addr); //checked

	//sign extending module
	sign_extender immediate_extender(inst_3, clk, extended_immediate); //checked

	//shift left by 2'er module
	doubleLeftShift immediate_shifter(extended_immediate, shifted_extended_immediate, 1, clk); //checked

	//operational register module
	//async_register register(read_1_addr, read_2_addr, write_addr, write_data, write_enable, read_1, read_2);
	regfile register(read_1, read_2, write_data, rs, rt, write_addr, write_enable, clk); //checked

	//alu source mux
	mux #(32) alu_src_mux(read_2, extended_immediate, alu_src, b); //checked 

	//alu module
	//alu ALU(a, b, alu_res, zero_flag);
	alu ALU(alu_res, carryout, zero_flag, overflow, read_1, b, alu_op); //checked

	//data memory module
	//data_memory data_mem(clk, mem_read_addr, mem_write_addr, mem_read_enable, mem_write_enable, mem_write_data_in, mem_read_data_out);
	datamemory data_memory(clk, alu_res, alu_res, mem_read_enable, mem_write_enable, read_2, mem_read); //checked

	//memory to register mux
	mux #(32) mem_to_reg_mux(alu_res, mem_read, mem_to_reg, normal_write_data); //checked

	//Optionally forces register to write PC+4 to whatever address
	//useful for jal operations
	mux #(32) jal_data_mux(normal_write_data, instruction_addr_plus4, jal_reg_override, write_data); //checked

endmodule
